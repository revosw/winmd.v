module metadata

pub struct Guid {
	data1 u32
	data2 u16
	data3 u16
	data4 [8]u8
}

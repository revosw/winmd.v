// module main

// #flag -lruntimeobject
// #flag -lrometadata

// fn C.RoInitialize(RoInitType) u32
// fn C.RoUninitialize()

// enum RoInitType {
// 	singlethreaded
// 	multithreaded
// }
